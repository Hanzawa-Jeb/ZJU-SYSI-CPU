`include "core_struct.vh"

module MaskGen(
    input CorePack::mem_op_enum mem_op,
    input CorePack::addr_t dmem_waddr,
    output CorePack::data_t dmem_wmask
);

  import CorePack::*;

  // Mask generation
  // fill your code

endmodule

