`ifdef VERILATE
    localparam FILE_PATH = "testcase.hex";
`else
    localparam FILE_PATH = ;// fill your testcase path
`endif